module OR_3 (in1,in2,in,out);
input in1,in2,in3;
output out;
    or U2(out,in1,in2,in3);
endmodule
